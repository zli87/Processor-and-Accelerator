
module MyDesign (
//---------------------------------------------------------------------------
//Control signals
          dut_run             ,
          dut_busy            ,
          reset_b             ,
          clk                 ,

//---------------------------------------------------------------------------
//input and output SRAM interface
          dut_sram_write_address  ,
          dut_sram_write_data     ,
          dut_sram_write_enable   ,
          dut_sram_read_address   ,
          sram_dut_read_data      ,
//---------------------------------------------------------------------------
//weights SRAM interface
          dut_wmem_read_address    ,
          wmem_dut_read_data
);

//---------------------------------------------------------------------------
//Control signals
input                 dut_run;
output  reg              dut_busy;
input                 reset_b;
input                 clk;

//---------------------------------------------------------------------------
//input and output SRAM interface
output   reg [11:0]       dut_sram_write_address;
output   reg [15:0]       dut_sram_write_data;
output   reg             dut_sram_write_enable;
output   reg [11:0]       dut_sram_read_address;
input    [15:0]       sram_dut_read_data;
//---------------------------------------------------------------------------
//weights SRAM interface
output   reg [11:0]       dut_wmem_read_address;
input    [15:0]       wmem_dut_read_data;

localparam  KERNEL_SIZE = 3;

localparam    S_IDLE = 3'b001;
localparam    S_FILL = 3'b010;
localparam    S_OUT = 3'b100;

reg [2:0] state_n;
reg [2:0] state_c;

reg [15:0] row0;
reg [15:0] row1;
reg [15:0] row2;
reg [9-1:0] weight;
reg [1:0] cnt_fill;
reg [1:0] dim; // 16: 10000,12: 01100, 10: 01010, compare index 4 and index 2
                //      10        01        00
reg [4:0] cnt_r;
reg [4:0] cnt_w;
reg flag_w;
wire flag_w_n ;
reg flag_last;
wire flag_last_n;
reg flag_r;
wire flag_r_n;
wire [1:0] read_offset;
wire [14-1:0] wdata;
wire [16-1:0] dut_sram_write_data_n;
wire [6-1:0] dut_sram_read_address_n;
wire [6-1:0] dut_sram_write_address_n;

always@(posedge clk or negedge reset_b)begin
    if(!reset_b)
        state_c<= 0;
    else
        state_c <= state_n;
end

always@(*) begin
    case(state_c)
        S_IDLE: if( dut_run ) state_n <= S_FILL;
                else state_n <= S_IDLE;
        S_FILL: if( &cnt_fill ) state_n <= S_OUT; //if(cnt_fill==2'd3)
                else state_n <= S_FILL;
        S_OUT:  if( flag_last ) state_n <= S_IDLE;
                else if( flag_w ) state_n <= S_FILL;
                else    state_n <= S_OUT;
        default: state_n <= S_IDLE;
    endcase
end
assign flag_last_n = ( flag_w_n )? (&row2[7:0]) : 1'b0; // row2 == 16'hff
always @ (posedge clk) begin
        flag_last <= flag_last_n;
end
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        cnt_fill <=0;
    else if( flag_w_n )
        cnt_fill <= 2'd3;
    else if(  state_c[1] )
        cnt_fill <= cnt_fill + 1;
    else if(!dut_busy)
        cnt_fill <= 0;
end
//==========================================================
// read weight
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        dut_wmem_read_address <= 12'd1;
    else
        dut_wmem_read_address <= 12'd1;
end
// weight == wmem_dut_read_data
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        weight <= 0;
    else
        weight <= wmem_dut_read_data[8:0];
end

//==========================================================
// read input

assign flag_r_n  = (dim[1])? (cnt_r==5'd15) // cnt_r == 15, max = 16
              : (dim[0])? (cnt_r==5'd11)   // cnt_r==11, max = 12 1011 1100
              :           (cnt_r==5'd09);  // cnt_r==9, max = 10
//assign flag_r_n  = (dim[1])? (cnt_r==5'd15)
//              : (dim[0])? (cnt_r==5'd11)
//              :           (cnt_r==5'd09);

always @ (posedge clk or negedge reset_b) begin
     if(!reset_b)
        flag_r <=0;
    else
        flag_r <= flag_r_n  ;
end

always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        cnt_r <=0;
    else if(  (state_c[0] & state_n[1]) | flag_r ) // dut_run
        cnt_r <= 0;
    else if(dut_busy)
        cnt_r <= cnt_r +1;
end

//assign read_offset = ((state_c[0] & state_n[1]) | (flag_r))? 2'd2 :
//                     ( dut_busy )? 2'd1 :
//                         2'd0;
assign read_offset[1] = ((state_c[0] & state_n[1]) | (flag_r));
assign read_offset[0] = ( dut_busy & (!flag_r)  );

assign  dut_sram_read_address_n = (flag_last)? 0 : dut_sram_read_address[5:0] + read_offset;
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        dut_sram_read_address <= 0;
    else
        //dut_sram_read_address <= {6'd0, !(flag_last)&(dut_sram_read_address[5]|dut_sram_read_address_n[5]),dut_sram_read_address_n[4:0]};
        dut_sram_read_address <= {6'd0, dut_sram_read_address_n};
end
always@(posedge clk or negedge reset_b)begin
    if(!reset_b)
        dim <= 0;
    else if( state_c[0] & state_n[1]  )
        dim <= {sram_dut_read_data[4], sram_dut_read_data[2]};
    else if( flag_w )
        dim <= {row1[4], row1[2]};
end
always@(posedge clk)begin
        row2 <= sram_dut_read_data;                     // input register
        row1 <= row2;                                   // pipeline register 1
        row0 <= row1;                                   // pipeline register 2
        dut_sram_write_data <= dut_sram_write_data_n ;  // output register
end
//==========================================================
// write output
assign flag_w_n = (dim[1])? (cnt_w==5'd13)
              : (dim[0])? (cnt_w==5'd9)
              :           (cnt_w==5'd7);
//assign flag_w_n = (dim[1])? (cnt_w==5'd13)
//              : (dim[0])? (cnt_w==5'd9)
//              :           (cnt_w==5'd7);
always @ (posedge clk) begin
    flag_w <= flag_w_n;
end
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        cnt_w <=0;
    else if(  (state_c[0] & state_n[1]) | (state_c[2] & state_n[1] ) ) // dut_run
        cnt_w <= 0;
    else if( dut_sram_write_enable )
        cnt_w <= cnt_w +1;
end

always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        dut_sram_write_enable <= 0;
    else if( flag_w_n | flag_w )
            dut_sram_write_enable <= 0;
    else if( state_c[2])
        dut_sram_write_enable <= 1;
end

assign dut_sram_write_address_n = dut_sram_write_address[4:0] + 1;
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        dut_sram_write_address <= 0;
    else if(state_c[2] & state_n[0])
        dut_sram_write_address <= 0;
    else if(dut_sram_write_enable)
        //dut_sram_write_address <= {6'd0, dut_sram_write_address_n[5] |dut_sram_write_address[5], dut_sram_write_address_n[4:0] };
        dut_sram_write_address <= {6'd0,dut_sram_write_address_n};
end
assign dut_sram_write_data_n =  (dim[1])? { 2'd0, wdata[14-1:0] }
                              : (dim[0])? { 6'd0, wdata[10-1:0] }
                              :           { 8'd0, wdata[8-1:0] };
genvar i;
wire [13:0] ans;
generate
    for(i=0;i<14;i=i+1)begin : pe
        PE inst( .w_i(weight), .A_i({ row2[i+2:i], row1[i+2:i], row0[i+2:i] }), .Z_o(wdata[i]) ); //, .ans(ans[i]) );
        //always @ (posedge clk) begin
        //        if(ans[i]!=wdata[i]) begin
        //            $display("xnor: %b, wdata[i]=%b, ans=%b",~(weight^{ row2[i+2:i], row1[i+2:i], row0[i+2:i] }),wdata[i],ans[i]);
        //            $finish;
        //        end
        //end
    end
endgenerate

// output busy signal
always @ (posedge clk or negedge reset_b) begin
    if(!reset_b)
        dut_busy <= 0;
    else if(flag_last_n)
        dut_busy <=0;
    else if(state_n[1])
        dut_busy <= 1;
end
endmodule

module PE(
    input [8:0] w_i,
    input [8:0] A_i,
    //output ans,
    output Z_o
);
wire [8:0] conv;
assign conv = ~(w_i^A_i);

//wire [3:0] sum; // max sum = 9 = 1001 > 4
//assign sum = conv[0] + conv[1] + conv[2] + conv[3] + conv[4] + conv[5] + conv[6] + conv[7] + conv[8];
// 0101 0110 0111 1000 1001
// sum[3] | (sum[2]&(sum[1]|sum[0]))
//assign ans = ( sum[3] | (sum[2]&(sum[1]|sum[0]) ) )? 1'b1 : 1'b0;

wire [1:0] sum1;
wire [1:0] sum2;
wire [1:0] sum3;
assign sum1 = conv[0]+conv[1]+conv[2];
assign sum2 = conv[3]+conv[4]+conv[5];
assign sum3 = conv[6]+conv[7]+conv[8];
// assume minimum of each sum
// 2,2,1|2  2,1|2,2  1|2,2,2
//3,1,1  1,3,1   1,1,3
// 3,2,?  2,3,? 3,?,2  2,?,3 ?,3,2  ?,2,3
/*
assign Z_o = (sum1[1]&sum2[1] & (sum3[1]|sum3[0])) | (sum1[1]& (sum2[1]|sum2[0]) &sum3[1]) | ((sum1[1]|sum1[0]) &sum2[1]&sum3[1]) |
        (sum1[1]&sum1[0] & sum2[0] & sum3[0]) | (sum1[0] & sum2[1]&sum2[0] & sum3[0]) | (sum1[0] & sum2[0] & sum3[1]&sum3[0]) |
        (sum1[1]&sum1[0] & sum2[1]) | (sum1[1] & sum2[1]&sum2[0]) |
        (sum1[1]&sum1[0] & sum3[1]) | (sum1[1] & sum3[1]&sum3[0]) |
        (sum2[1]&sum2[0] & sum3[1]) | (sum2[1] & sum3[1]&sum3[0]);
*/
assign Z_o = ( (sum1[1]|sum2[1]|sum3[1]) &sum1[0] & sum2[0] & sum3[0]) |
        (sum1[1]&sum2[1] & ((sum1[0]|sum2[0]|sum3[1]|sum3[0])) ) |
        (sum1[1]&sum3[1] & ((sum1[0]|sum3[0]|sum2[1]|sum2[0])) ) |
        (sum2[1]&sum3[1] & ((sum2[0]|sum3[0]|sum1[1]|sum1[0])) );

endmodule
